module hdmi_config_queue(

);

endmodule
